module test1(
	input wire clk,
	output wire clk1
);

assign clk1 = clk;

endmodule

